module initializing